library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity test_buff is
end entity test_buff;


architecture testing_buff of test_buff is


component Buffer_Module is
port (

	clk, reset: in std_logic;
	shift_enable : in std_logic;
	data_in : in std_logic_vector(7 downto 0);
	
	px1, px2, px3, px4, px5, px6, px7, px8, px9 : out std_logic_vector(7 downto 0)
		
);
end component Buffer_Module;



signal clk_s,enable_s, reset_s : std_logic := '0';

signal pix_in : std_logic_vector(7 downto 0) := (others => '0');

signal p1, p2, p3, p4, p5, p6, p7, p8, p9 : std_logic_vector(7 downto 0) := (others => '0');

--signal kern_sel_s : std_logic_vector(2 downto 0) := (others => '0');

--signal im_width : std_logic_vector(10 downto 0) := (others => '0');
--signal im_height : std_logic_vector(9 downto 0) := (others => '0');




begin

buffer_mod : Buffer_Module port map (

	clk => clk_s,
	reset => reset_s,
	shift_enable => enable_s,
	data_in => pix_in,
	px1 => p1,
	px2 => p2,
	px3 => p3,
	px4 => p4,
	px5 => p5,
	px6 => p6,
	px7 => p7,
	px8 => p8,
	px9 => p9

);




	timing : process
	begin
	
		wait for 2 ns;
		clk_s <= '1';
		wait for 2 ns;
		clk_s <= '0';

	end process;
	
	data : process
	begin
	
	--reset_s <= '1', '0' after 2 ns;	
	
	enable_s <= '0', '1' after 4 ns, '0' after 39 ns , '1' after 54 ns, '0' after 82 ns;
	
	pix_in <= x"00" after 4 ns, 
					x"00" after 8 ns, 
					x"FF" after 12 ns, 
					x"00" after 16 ns, 
					x"00" after 20 ns, 
					x"00" after 24 ns, 
					x"FF" after 28 ns, 
					x"FF" after 32 ns, 
					x"00" after 36 ns, 
					x"00" after 40 ns, 
					x"00" after 44 ns, 
					x"00" after 48 ns, 
					x"FF" after 52 ns, 
					x"00" after 56 ns, 
					x"00" after 60 ns, 
					x"00" after 64 ns, 
					x"00" after 68 ns, 
					x"FF" after 72 ns, 
					x"00" after 76 ns, 
					x"00" after 80 ns, 
					x"FF" after 84 ns, 
					x"FF" after 88 ns, 
					x"FF" after 92 ns, 
					x"FF" after 96 ns, 
					x"FF" after 100 ns;	
	wait;
	
	end process;
	

end architecture testing_buff;